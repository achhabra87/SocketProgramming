-- Copyright (C) 1991-2007 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 7.2 Build 151 09/26/2007 SJ Full Version
-- Created on Sun Feb 12 22:52:16 2012

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SM1 IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        input1 : IN STD_LOGIC := '0';
        input2 : IN STD_LOGIC := '0';
        output1 : OUT STD_LOGIC
    );
END SM1;

ARCHITECTURE BEHAVIOR OF SM1 IS
    TYPE type_fstate IS (state2,state3,state1);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
    SIGNAL reg_output1 : STD_LOGIC := '0';
BEGIN
    PROCESS (clock,reg_fstate,reg_output1)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
            output1 <= reg_output1;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,input1,input2)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state1;
            reg_output1 <= '0';
        ELSE
            CASE fstate IS
                WHEN state2 =>
                    IF (((input1 = '1') AND NOT((input2 = '1')))) THEN
                        reg_fstate <= state3;
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    reg_output1 <= '0';
                WHEN state3 =>
                    IF (((input1 = '1') OR (input2 = '1'))) THEN
                        reg_fstate <= state1;
                    ELSE
                        reg_fstate <= state3;
                    END IF;

                    reg_output1 <= '1';
                WHEN state1 =>
                    IF (((input1 = '1') AND (input2 = '1'))) THEN
                        reg_fstate <= state2;
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    reg_output1 <= '1';
                WHEN OTHERS => 
                    reg_output1 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
